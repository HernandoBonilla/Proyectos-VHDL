-- Library and packages 
library	IEEE;
use IEEE.std_logic_1164.all;

-- Entity (empty)
entity mux8way_test is	
end entity;

-- Architecture (test process)
architecture arch_test of mux8way_test is

	-- Component declaration
	component mux8way
		port(
			a	:	in 	std_logic;
			b	:	in		std_logic;
			c 	: 	in 	std_logic;
			d	: 	in 	std_logic;
			e	: 	in 	std_logic;
			f	:	in		std_logic;
			g	:	in		std_logic;
			h	:	in		std_logic;
			s1 :	in 	std_logic;
			s2 : 	in 	std_logic;
			s3 : 	in 	std_logic;
			o	:	out	std_logic
		);
	end component;
	
	-- Signal declaration
	signal a_test		: std_logic := '0';
	signal b_test		: std_logic := '0';
	signal c_test		: std_logic := '0';
	signal d_test		: std_logic := '0';
	signal e_test		: std_logic := '0';
	signal f_test		: std_logic := '0';
	signal g_test		: std_logic := '0';
	signal h_test		: std_logic := '0';
	signal s1_test	   : std_logic := '0';
	signal s2_test		: std_logic := '0';
	signal s3_test 	: std_logic := '0';
	signal o_test		: std_logic;
	
	begin
	
	-- DUT instantiation
	dut1	: mux8way 
		port map (
			a 		=> a_test,
			b 		=> b_test,
			c		=> c_test,
			d 		=> d_test,
			e 		=> e_test,
			f 		=> f_test,
			g		=> g_test,
			h 		=> h_test,
			s1		=> s1_test,
			s2 	=> s2_test,
			s3		=> s3_test,
			o 		=> o_test
		);

	-- Stimulus generation
	Stimulus	: process
	begin
	  
	   report "Start of the test of mux4way"	  
		severity note;
		
		a_test 	<= '0';
		b_test 	<= '0';
		c_test 	<= '0';
		d_test   <= '1';
		e_test 	<= '0';
		f_test 	<= '0';
		g_test 	<= '0';
		h_test   <= '1';
		s1_test  <= '0';
		s2_test	<= '0';
		s3_test  <= '0';
		wait for 1 ns;
		assert o_test = '1'
		  report "Failure for {a,b,c,d,e,f,g,h,s1,s2,s3} = {0,0,0,0,0,0,0,1,0,0,0}"
		  severity failure;
		  
		a_test 	<= '0';
		b_test 	<= '0';
		c_test 	<= '0';
		d_test   <= '0';
		e_test 	<= '0';
		f_test 	<= '0';
		g_test 	<= '1';
		h_test   <= '0';
		s1_test  <= '0';
		s2_test	<= '0';
		s3_test  <= '1';
		wait for 1 ns;
		assert o_test = '1'
		  report "Failure for {a,b,c,d,e,f,g,h,s1,s2,s3} = {0,0,0,0,0,0,1,0,0,0,1}"
		  severity failure;
		
		a_test 	<= '0';
		b_test 	<= '0';
		c_test 	<= '0';
		d_test   <= '0';
		e_test 	<= '0';
		f_test 	<= '1';
		g_test 	<= '0';
		h_test   <= '0';
		s1_test  <= '0';
		s2_test	<= '1';
		s3_test  <= '0';
		wait for 1 ns;
		assert o_test = '1'
		  report "Failure for {a,b,c,d,e,f,g,h,s1,s2,s3} = {0,0,0,0,0,1,0,0,0,1,0}"
		  severity failure;	  

		a_test 	<= '0';
		b_test 	<= '0';
		c_test 	<= '0';
		d_test   <= '0';
		e_test 	<= '1';
		f_test 	<= '0';
		g_test 	<= '0';
		h_test   <= '0';
		s1_test  <= '0';
		s2_test	<= '1';
		s3_test  <= '1';
		wait for 1 ns;
		assert o_test = '1'
		  report "Failure for {a,b,c,d,e,f,g,h,s1,s2,s3} = {0,0,0,0,1,0,0,0,0,1,1}"
		  severity failure;
		
		a_test 	<= '0';
		b_test 	<= '0';
		c_test 	<= '0';
		d_test   <= '1';
		e_test 	<= '0';
		f_test 	<= '0';
		g_test 	<= '0';
		h_test   <= '0';
		s1_test  <= '1';
		s2_test	<= '0';
		s3_test  <= '0';
		wait for 1 ns;
		assert o_test = '1'
		  report "Failure for {a,b,c,d,e,f,g,h,s1,s2,s3} = {0,0,0,1,0,0,0,0,1,0,0}"
		  severity failure;
		  
		a_test 	<= '0';
		b_test 	<= '0';
		c_test 	<= '1';
		d_test   <= '0';
		e_test 	<= '0';
		f_test 	<= '0';
		g_test 	<= '0';
		h_test   <= '0';
		s1_test  <= '1';
		s2_test	<= '0';
		s3_test  <= '1';
		wait for 1 ns;
		assert o_test = '1'
		  report "Failure for {a,b,c,d,e,f,g,h,s1,s2,s3} = {0,0,1,0,0,0,0,0,1,0,1}"
		  severity failure;
		  
		a_test 	<= '0';
		b_test 	<= '1';
		c_test 	<= '0';
		d_test   <= '0';
		e_test 	<= '0';
		f_test 	<= '0';
		g_test 	<= '0';
		h_test   <= '0';
		s1_test  <= '1';
		s2_test	<= '1';
		s3_test  <= '0';
		wait for 1 ns;
		assert o_test = '1'
		  report "Failure for {a,b,c,d,e,f,g,h,s1,s2,s3} = {0,1,0,0,0,0,0,0,1,1,0}"
		  severity failure;
		  
		a_test 	<= '1';
		b_test 	<= '0';
		c_test 	<= '0';
		d_test   <= '0';
		e_test 	<= '0';
		f_test 	<= '0';
		g_test 	<= '0';
		h_test   <= '0';
		s1_test  <= '1';
		s2_test	<= '1';
		s3_test  <= '1';
		wait for 1 ns;
		assert o_test = '1'
		  report "Failure for {a,b,c,d,e,f,g,h,s1,s2,s3} = {1,0,0,0,0,0,0,0,1,1,1}"
		  severity failure;
		  
		  
		a_test 	<= '0';
		b_test 	<= '1';
		c_test 	<= '0';
		d_test   <= '1';
		e_test 	<= '1';
		f_test 	<= '1';
		g_test 	<= '1';
		h_test   <= '0';
		s1_test  <= '1';
		s2_test	<= '1';
		s3_test  <= '1';
		wait for 1 ns;
		assert o_test = '0'
		  report "Failure for {a,b,c,d,e,f,g,h,s1,s2,s3} = {0,1,0,1,1,1,1,0,1,1,1}"
		  severity failure;
		  
		report "Test successful"
		severity note;
		wait;
		
	end process;

end architecture;